`include "4bit_adder.v"

module  adder_tb;
    reg[3;0]    x,y;
    wire[3:0]   s;
    wire        c_out;
    

