//--------------------------------------//
// Encoder con prioridad de 4 inputs    //
// Nombre del archivo: encoder_x4.v     //
// Electronica III - Grupo 4            //
// -------------------------------------//

module encoder_x4(z1, z2, y, x);
    
    // Inputs-Outputs
    input[3:0]  x;
    output      z1, z2, y;
    wire        z1, z2, y;

    // Descripción de nodos internos
    wire        net1, net2;
endmodule