module two_complement_adder();


// Sumador con entrada de control M.
// Si M = 1, hace XOR(1;y_i) y obtengo el Complemento a 1 de Y
// en las entradas.
// Pongo el C_-1 en M = 1 para obtener el complemento a 2 de Y.
// Sumo X + C_2(Y).

// Si obtengo Carry (salida negada) significa que X<Y, de lo contrario X>=Y
// Hago el circuito para todos los flags (S,Z,V,C)


endmodule